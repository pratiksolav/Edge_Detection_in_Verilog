module test_just_2(bus,bus_con,clk,reset,strobe_data,strobe_mode);
inout [7:0]bus;
input strobe_data,strobe_mode,bus_con,reset,clk;
wire [7:0]bus_1;
reg [7:0]bus_2;

reg [7:0]r1[121:0];
reg [7:0]r2[121:0];
reg [7:0]r3[121:0];

reg [6:0]Windex,Rindex,i;
reg write,read;
assign bus=(bus_con)?bus_2:8'dz;
assign bus_1=(!bus_con)?bus:8'dz;

wire [7:0]edges[119:0];
sobel_edge A0(r1[0],r1[1],r1[2],r2[0],r2[2],r3[0],r3[1],r3[2],edges[0]);
sobel_edge A1(r1[1],r1[2],r1[3],r2[1],r2[3],r3[1],r3[2],r3[3],edges[1]);
sobel_edge A2(r1[2],r1[3],r1[4],r2[2],r2[4],r3[2],r3[3],r3[4],edges[2]);
sobel_edge A3(r1[3],r1[4],r1[5],r2[3],r2[5],r3[3],r3[4],r3[5],edges[3]);
sobel_edge A4(r1[4],r1[5],r1[6],r2[4],r2[6],r3[4],r3[5],r3[6],edges[4]);
sobel_edge A5(r1[5],r1[6],r1[7],r2[5],r2[7],r3[5],r3[6],r3[7],edges[5]);
sobel_edge A6(r1[6],r1[7],r1[8],r2[6],r2[8],r3[6],r3[7],r3[8],edges[6]);
sobel_edge A7(r1[7],r1[8],r1[9],r2[7],r2[9],r3[7],r3[8],r3[9],edges[7]);
sobel_edge A8(r1[8],r1[9],r1[10],r2[8],r2[10],r3[8],r3[9],r3[10],edges[8]);
sobel_edge A9(r1[9],r1[10],r1[11],r2[9],r2[11],r3[9],r3[10],r3[11],edges[9]);
sobel_edge A10(r1[10],r1[11],r1[12],r2[10],r2[12],r3[10],r3[11],r3[12],edges[10]);
sobel_edge A11(r1[11],r1[12],r1[13],r2[11],r2[13],r3[11],r3[12],r3[13],edges[11]);
sobel_edge A12(r1[12],r1[13],r1[14],r2[12],r2[14],r3[12],r3[13],r3[14],edges[12]);
sobel_edge A13(r1[13],r1[14],r1[15],r2[13],r2[15],r3[13],r3[14],r3[15],edges[13]);
sobel_edge A14(r1[14],r1[15],r1[16],r2[14],r2[16],r3[14],r3[15],r3[16],edges[14]);
sobel_edge A15(r1[15],r1[16],r1[17],r2[15],r2[17],r3[15],r3[16],r3[17],edges[15]);
sobel_edge A16(r1[16],r1[17],r1[18],r2[16],r2[18],r3[16],r3[17],r3[18],edges[16]);
sobel_edge A17(r1[17],r1[18],r1[19],r2[17],r2[19],r3[17],r3[18],r3[19],edges[17]);
sobel_edge A18(r1[18],r1[19],r1[20],r2[18],r2[20],r3[18],r3[19],r3[20],edges[18]);
sobel_edge A19(r1[19],r1[20],r1[21],r2[19],r2[21],r3[19],r3[20],r3[21],edges[19]);
sobel_edge A20(r1[20],r1[21],r1[22],r2[20],r2[22],r3[20],r3[21],r3[22],edges[20]);
sobel_edge A21(r1[21],r1[22],r1[23],r2[21],r2[23],r3[21],r3[22],r3[23],edges[21]);
sobel_edge A22(r1[22],r1[23],r1[24],r2[22],r2[24],r3[22],r3[23],r3[24],edges[22]);
sobel_edge A23(r1[23],r1[24],r1[25],r2[23],r2[25],r3[23],r3[24],r3[25],edges[23]);
sobel_edge A24(r1[24],r1[25],r1[26],r2[24],r2[26],r3[24],r3[25],r3[26],edges[24]);
sobel_edge A25(r1[25],r1[26],r1[27],r2[25],r2[27],r3[25],r3[26],r3[27],edges[25]);
sobel_edge A26(r1[26],r1[27],r1[28],r2[26],r2[28],r3[26],r3[27],r3[28],edges[26]);
sobel_edge A27(r1[27],r1[28],r1[29],r2[27],r2[29],r3[27],r3[28],r3[29],edges[27]);
sobel_edge A28(r1[28],r1[29],r1[30],r2[28],r2[30],r3[28],r3[29],r3[30],edges[28]);
sobel_edge A29(r1[29],r1[30],r1[31],r2[29],r2[31],r3[29],r3[30],r3[31],edges[29]);
sobel_edge A30(r1[30],r1[31],r1[32],r2[30],r2[32],r3[30],r3[31],r3[32],edges[30]);
sobel_edge A31(r1[31],r1[32],r1[33],r2[31],r2[33],r3[31],r3[32],r3[33],edges[31]);
sobel_edge A32(r1[32],r1[33],r1[34],r2[32],r2[34],r3[32],r3[33],r3[34],edges[32]);
sobel_edge A33(r1[33],r1[34],r1[35],r2[33],r2[35],r3[33],r3[34],r3[35],edges[33]);
sobel_edge A34(r1[34],r1[35],r1[36],r2[34],r2[36],r3[34],r3[35],r3[36],edges[34]);
sobel_edge A35(r1[35],r1[36],r1[37],r2[35],r2[37],r3[35],r3[36],r3[37],edges[35]);
sobel_edge A36(r1[36],r1[37],r1[38],r2[36],r2[38],r3[36],r3[37],r3[38],edges[36]);
sobel_edge A37(r1[37],r1[38],r1[39],r2[37],r2[39],r3[37],r3[38],r3[39],edges[37]);
sobel_edge A38(r1[38],r1[39],r1[40],r2[38],r2[40],r3[38],r3[39],r3[40],edges[38]);
sobel_edge A39(r1[39],r1[40],r1[41],r2[39],r2[41],r3[39],r3[40],r3[41],edges[39]);
sobel_edge A40(r1[40],r1[41],r1[42],r2[40],r2[42],r3[40],r3[41],r3[42],edges[40]);
sobel_edge A41(r1[41],r1[42],r1[43],r2[41],r2[43],r3[41],r3[42],r3[43],edges[41]);
sobel_edge A42(r1[42],r1[43],r1[44],r2[42],r2[44],r3[42],r3[43],r3[44],edges[42]);
sobel_edge A43(r1[43],r1[44],r1[45],r2[43],r2[45],r3[43],r3[44],r3[45],edges[43]);
sobel_edge A44(r1[44],r1[45],r1[46],r2[44],r2[46],r3[44],r3[45],r3[46],edges[44]);
sobel_edge A45(r1[45],r1[46],r1[47],r2[45],r2[47],r3[45],r3[46],r3[47],edges[45]);
sobel_edge A46(r1[46],r1[47],r1[48],r2[46],r2[48],r3[46],r3[47],r3[48],edges[46]);
sobel_edge A47(r1[47],r1[48],r1[49],r2[47],r2[49],r3[47],r3[48],r3[49],edges[47]);
sobel_edge A48(r1[48],r1[49],r1[50],r2[48],r2[50],r3[48],r3[49],r3[50],edges[48]);
sobel_edge A49(r1[49],r1[50],r1[51],r2[49],r2[51],r3[49],r3[50],r3[51],edges[49]);
sobel_edge A50(r1[50],r1[51],r1[52],r2[50],r2[52],r3[50],r3[51],r3[52],edges[50]);
sobel_edge A51(r1[51],r1[52],r1[53],r2[51],r2[53],r3[51],r3[52],r3[53],edges[51]);
sobel_edge A52(r1[52],r1[53],r1[54],r2[52],r2[54],r3[52],r3[53],r3[54],edges[52]);
sobel_edge A53(r1[53],r1[54],r1[55],r2[53],r2[55],r3[53],r3[54],r3[55],edges[53]);
sobel_edge A54(r1[54],r1[55],r1[56],r2[54],r2[56],r3[54],r3[55],r3[56],edges[54]);
sobel_edge A55(r1[55],r1[56],r1[57],r2[55],r2[57],r3[55],r3[56],r3[57],edges[55]);
sobel_edge A56(r1[56],r1[57],r1[58],r2[56],r2[58],r3[56],r3[57],r3[58],edges[56]);
sobel_edge A57(r1[57],r1[58],r1[59],r2[57],r2[59],r3[57],r3[58],r3[59],edges[57]);
sobel_edge A58(r1[58],r1[59],r1[60],r2[58],r2[60],r3[58],r3[59],r3[60],edges[58]);
sobel_edge A59(r1[59],r1[60],r1[61],r2[59],r2[61],r3[59],r3[60],r3[61],edges[59]);
sobel_edge A60(r1[60],r1[61],r1[62],r2[60],r2[62],r3[60],r3[61],r3[62],edges[60]);
sobel_edge A61(r1[61],r1[62],r1[63],r2[61],r2[63],r3[61],r3[62],r3[63],edges[61]);
sobel_edge A62(r1[62],r1[63],r1[64],r2[62],r2[64],r3[62],r3[63],r3[64],edges[62]);
sobel_edge A63(r1[63],r1[64],r1[65],r2[63],r2[65],r3[63],r3[64],r3[65],edges[63]);
sobel_edge A64(r1[64],r1[65],r1[66],r2[64],r2[66],r3[64],r3[65],r3[66],edges[64]);
sobel_edge A65(r1[65],r1[66],r1[67],r2[65],r2[67],r3[65],r3[66],r3[67],edges[65]);
sobel_edge A66(r1[66],r1[67],r1[68],r2[66],r2[68],r3[66],r3[67],r3[68],edges[66]);
sobel_edge A67(r1[67],r1[68],r1[69],r2[67],r2[69],r3[67],r3[68],r3[69],edges[67]);
sobel_edge A68(r1[68],r1[69],r1[70],r2[68],r2[70],r3[68],r3[69],r3[70],edges[68]);
sobel_edge A69(r1[69],r1[70],r1[71],r2[69],r2[71],r3[69],r3[70],r3[71],edges[69]);
sobel_edge A70(r1[70],r1[71],r1[72],r2[70],r2[72],r3[70],r3[71],r3[72],edges[70]);
sobel_edge A71(r1[71],r1[72],r1[73],r2[71],r2[73],r3[71],r3[72],r3[73],edges[71]);
sobel_edge A72(r1[72],r1[73],r1[74],r2[72],r2[74],r3[72],r3[73],r3[74],edges[72]);
sobel_edge A73(r1[73],r1[74],r1[75],r2[73],r2[75],r3[73],r3[74],r3[75],edges[73]);
sobel_edge A74(r1[74],r1[75],r1[76],r2[74],r2[76],r3[74],r3[75],r3[76],edges[74]);
sobel_edge A75(r1[75],r1[76],r1[77],r2[75],r2[77],r3[75],r3[76],r3[77],edges[75]);
sobel_edge A76(r1[76],r1[77],r1[78],r2[76],r2[78],r3[76],r3[77],r3[78],edges[76]);
sobel_edge A77(r1[77],r1[78],r1[79],r2[77],r2[79],r3[77],r3[78],r3[79],edges[77]);
sobel_edge A78(r1[78],r1[79],r1[80],r2[78],r2[80],r3[78],r3[79],r3[80],edges[78]);
sobel_edge A79(r1[79],r1[80],r1[81],r2[79],r2[81],r3[79],r3[80],r3[81],edges[79]);
sobel_edge A80(r1[80],r1[81],r1[82],r2[80],r2[82],r3[80],r3[81],r3[82],edges[80]);
sobel_edge A81(r1[81],r1[82],r1[83],r2[81],r2[83],r3[81],r3[82],r3[83],edges[81]);
sobel_edge A82(r1[82],r1[83],r1[84],r2[82],r2[84],r3[82],r3[83],r3[84],edges[82]);
sobel_edge A83(r1[83],r1[84],r1[85],r2[83],r2[85],r3[83],r3[84],r3[85],edges[83]);
sobel_edge A84(r1[84],r1[85],r1[86],r2[84],r2[86],r3[84],r3[85],r3[86],edges[84]);
sobel_edge A85(r1[85],r1[86],r1[87],r2[85],r2[87],r3[85],r3[86],r3[87],edges[85]);
sobel_edge A86(r1[86],r1[87],r1[88],r2[86],r2[88],r3[86],r3[87],r3[88],edges[86]);
sobel_edge A87(r1[87],r1[88],r1[89],r2[87],r2[89],r3[87],r3[88],r3[89],edges[87]);
sobel_edge A88(r1[88],r1[89],r1[90],r2[88],r2[90],r3[88],r3[89],r3[90],edges[88]);
sobel_edge A89(r1[89],r1[90],r1[91],r2[89],r2[91],r3[89],r3[90],r3[91],edges[89]);
sobel_edge A90(r1[90],r1[91],r1[92],r2[90],r2[92],r3[90],r3[91],r3[92],edges[90]);
sobel_edge A91(r1[91],r1[92],r1[93],r2[91],r2[93],r3[91],r3[92],r3[93],edges[91]);
sobel_edge A92(r1[92],r1[93],r1[94],r2[92],r2[94],r3[92],r3[93],r3[94],edges[92]);
sobel_edge A93(r1[93],r1[94],r1[95],r2[93],r2[95],r3[93],r3[94],r3[95],edges[93]);
sobel_edge A94(r1[94],r1[95],r1[96],r2[94],r2[96],r3[94],r3[95],r3[96],edges[94]);
sobel_edge A95(r1[95],r1[96],r1[97],r2[95],r2[97],r3[95],r3[96],r3[97],edges[95]);
sobel_edge A96(r1[96],r1[97],r1[98],r2[96],r2[98],r3[96],r3[97],r3[98],edges[96]);
sobel_edge A97(r1[97],r1[98],r1[99],r2[97],r2[99],r3[97],r3[98],r3[99],edges[97]);
sobel_edge A98(r1[98],r1[99],r1[100],r2[98],r2[100],r3[98],r3[99],r3[100],edges[98]);
sobel_edge A99(r1[99],r1[100],r1[101],r2[99],r2[101],r3[99],r3[100],r3[101],edges[99]);
sobel_edge A100(r1[100],r1[101],r1[102],r2[100],r2[102],r3[100],r3[101],r3[102],edges[100]);
sobel_edge A101(r1[101],r1[102],r1[103],r2[101],r2[103],r3[101],r3[102],r3[103],edges[101]);
sobel_edge A102(r1[102],r1[103],r1[104],r2[102],r2[104],r3[102],r3[103],r3[104],edges[102]);
sobel_edge A103(r1[103],r1[104],r1[105],r2[103],r2[105],r3[103],r3[104],r3[105],edges[103]);
sobel_edge A104(r1[104],r1[105],r1[106],r2[104],r2[106],r3[104],r3[105],r3[106],edges[104]);
sobel_edge A105(r1[105],r1[106],r1[107],r2[105],r2[107],r3[105],r3[106],r3[107],edges[105]);
sobel_edge A106(r1[106],r1[107],r1[108],r2[106],r2[108],r3[106],r3[107],r3[108],edges[106]);
sobel_edge A107(r1[107],r1[108],r1[109],r2[107],r2[109],r3[107],r3[108],r3[109],edges[107]);
sobel_edge A108(r1[108],r1[109],r1[110],r2[108],r2[110],r3[108],r3[109],r3[110],edges[108]);
sobel_edge A109(r1[109],r1[110],r1[111],r2[109],r2[111],r3[109],r3[110],r3[111],edges[109]);
sobel_edge A110(r1[110],r1[111],r1[112],r2[110],r2[112],r3[110],r3[111],r3[112],edges[110]);
sobel_edge A111(r1[111],r1[112],r1[113],r2[111],r2[113],r3[111],r3[112],r3[113],edges[111]);
sobel_edge A112(r1[112],r1[113],r1[114],r2[112],r2[114],r3[112],r3[113],r3[114],edges[112]);
sobel_edge A113(r1[113],r1[114],r1[115],r2[113],r2[115],r3[113],r3[114],r3[115],edges[113]);
sobel_edge A114(r1[114],r1[115],r1[116],r2[114],r2[116],r3[114],r3[115],r3[116],edges[114]);
sobel_edge A115(r1[115],r1[116],r1[117],r2[115],r2[117],r3[115],r3[116],r3[117],edges[115]);
sobel_edge A116(r1[116],r1[117],r1[118],r2[116],r2[118],r3[116],r3[117],r3[118],edges[116]);
sobel_edge A117(r1[117],r1[118],r1[119],r2[117],r2[119],r3[117],r3[118],r3[119],edges[117]);
sobel_edge A118(r1[118],r1[119],r1[120],r2[118],r2[120],r3[118],r3[119],r3[120],edges[118]);
sobel_edge A119(r1[119],r1[120],r1[121],r2[119],r2[121],r3[119],r3[120],r3[121],edges[119]);

always@(posedge clk,negedge reset)
begin
if(!reset)
begin
Windex<=7'b0;Rindex<=7'b0;read<=1'b0;write<=1'b0;
for(i=0;i<122;i=i+1)
begin
r1[i]<=8'b0;
r2[i]<=8'b0;
end
bus_2<=8'hff;
end
else if(!strobe_data &!bus_con&!write)
begin
r3[Windex]<=bus_1;
Windex<=Windex+1;
write<=1'b0;
end
else if(!strobe_data & bus_con & !read)
begin
case(Rindex+1)
  1:bus_2<=edges[0];  
 2:bus_2<=edges[1];  
 3:bus_2<=edges[2];  
 4:bus_2<=edges[3];  
 5:bus_2<=edges[4];  
 6:bus_2<=edges[5];  
 7:bus_2<=edges[6];  
 8:bus_2<=edges[7];  
 9:bus_2<=edges[8];  
 10:bus_2<=edges[9];  
 11:bus_2<=edges[10];  
 12:bus_2<=edges[11];  
 13:bus_2<=edges[12];  
 14:bus_2<=edges[13];  
 15:bus_2<=edges[14];  
 16:bus_2<=edges[15];  
 17:bus_2<=edges[16];  
 18:bus_2<=edges[17];  
 19:bus_2<=edges[18];  
 20:bus_2<=edges[19];  
 21:bus_2<=edges[20];  
 22:bus_2<=edges[21];  
 23:bus_2<=edges[22];  
 24:bus_2<=edges[23];  
 25:bus_2<=edges[24];  
 26:bus_2<=edges[25];  
 27:bus_2<=edges[26];  
 28:bus_2<=edges[27];  
 29:bus_2<=edges[28];  
 30:bus_2<=edges[29];  
 31:bus_2<=edges[30];  
 32:bus_2<=edges[31];  
 33:bus_2<=edges[32];  
 34:bus_2<=edges[33];  
 35:bus_2<=edges[34];  
 36:bus_2<=edges[35];  
 37:bus_2<=edges[36];  
 38:bus_2<=edges[37];  
 39:bus_2<=edges[38];  
 40:bus_2<=edges[39];  
 41:bus_2<=edges[40];  
 42:bus_2<=edges[41];  
 43:bus_2<=edges[42];  
 44:bus_2<=edges[43];  
 45:bus_2<=edges[44];  
 46:bus_2<=edges[45];  
 47:bus_2<=edges[46];  
 48:bus_2<=edges[47];  
 49:bus_2<=edges[48];  
 50:bus_2<=edges[49];  
 51:bus_2<=edges[50];  
 52:bus_2<=edges[51];  
 53:bus_2<=edges[52];  
 54:bus_2<=edges[53];  
 55:bus_2<=edges[54];  
 56:bus_2<=edges[55];  
 57:bus_2<=edges[56];  
 58:bus_2<=edges[57];  
 59:bus_2<=edges[58];  
 60:bus_2<=edges[59];  
 61:bus_2<=edges[60];  
 62:bus_2<=edges[61];  
 63:bus_2<=edges[62];  
 64:bus_2<=edges[63];  
 65:bus_2<=edges[64];  
 66:bus_2<=edges[65];  
 67:bus_2<=edges[66];  
 68:bus_2<=edges[67];  
 69:bus_2<=edges[68];  
 70:bus_2<=edges[69];  
 71:bus_2<=edges[70];  
 72:bus_2<=edges[71];  
 73:bus_2<=edges[72];  
 74:bus_2<=edges[73];  
 75:bus_2<=edges[74];  
 76:bus_2<=edges[75];  
 77:bus_2<=edges[76];  
 78:bus_2<=edges[77];  
 79:bus_2<=edges[78];  
 80:bus_2<=edges[79];  
 81:bus_2<=edges[80];  
 82:bus_2<=edges[81];  
 83:bus_2<=edges[82];  
 84:bus_2<=edges[83];  
 85:bus_2<=edges[84];  
 86:bus_2<=edges[85];  
 87:bus_2<=edges[86];  
 88:bus_2<=edges[87];  
 89:bus_2<=edges[88];  
 90:bus_2<=edges[89];  
 91:bus_2<=edges[90];  
 92:bus_2<=edges[91];  
 93:bus_2<=edges[92];  
 94:bus_2<=edges[93];  
 95:bus_2<=edges[94];  
 96:bus_2<=edges[95];  
 97:bus_2<=edges[96];  
 98:bus_2<=edges[97];  
 99:bus_2<=edges[98];  
 100:bus_2<=edges[99];  
 101:bus_2<=edges[100];  
 102:bus_2<=edges[101];  
 103:bus_2<=edges[102];  
 104:bus_2<=edges[103];  
 105:bus_2<=edges[104];  
 106:bus_2<=edges[105];  
 107:bus_2<=edges[106];  
 108:bus_2<=edges[107];  
 109:bus_2<=edges[108];  
 110:bus_2<=edges[109];  
 111:bus_2<=edges[110];  
 112:bus_2<=edges[111];  
 113:bus_2<=edges[112];  
 114:bus_2<=edges[113];  
 115:bus_2<=edges[114];  
 116:bus_2<=edges[115];  
 117:bus_2<=edges[116];  
 118:bus_2<=edges[117];  
 119:bus_2<=edges[118];  
 120:bus_2<=edges[119];  
  default:bus_2<=8'b0;
endcase
Rindex<=Rindex+1;
read<=1'b0;
end
else if(!strobe_mode & !bus_con & !write)
begin
for(i=0;i<122;i=i+1)
begin
r1[i]<=r2[i];
r2[i]<=r3[i];
end
Windex<=7'b0;
Rindex<=7'b0;
write<=1'b0;
bus_2<=8'b0;
end
end
endmodule
module sobel_edge(pix0,pix1,pix2,pix3,pix5,pix6,pix7,pix8,edges);
input  [7:0]pix0,pix1,pix2,pix3,pix5,pix6,pix7,pix8;	
output [7:0]edges;				
wire signed [10:0]x,y;  					 
wire signed [10:0]mod_x,mod_y;
wire [10:0]sum;
assign x=((pix2-pix0)+((pix5-pix3)<<1)+(pix8-pix6)); 
assign y=((pix0-pix6)+((pix1-pix7)<<1)+(pix2-pix8));
assign mod_x=(x[10]?~x+1:x);	 
assign mod_y=(y[10]?~y+1:y); 
assign sum = (mod_x+mod_y);			
assign edges=(sum[10:8])?8'hff:sum[7:0];	
endmodule
